LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ji IS
PORT(
SW:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
LED:OUT STD_LOGIC);
END;
ARCHITECTURE A OF ji IS
BEGIN
LED <= SW(0) XOR SW(1) XOR SW(2) XOR SW(3);
END;