LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY zcc IS
PORT(
clk:IN STD_LOGIC;
seg:OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
c:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END zcc;
ARCHITECTURE A OF zcc IS
SIGNAL S:INTEGER RANGE 0 TO 7;

BEGIN
PROCESS(clk,S)
BEGIN
IF clk'EVENT AND clk='1'THEN
IF S=7 THEN
  S<=0;
ELSE S<=S+1;
END IF;
END IF;
END PROCESS;



PROCESS(S)
BEGIN
case S IS
WHEN 0=>c<="01111111";seg<="0110000";--1
WHEN 1=>c<="10111111";seg<="1011111";--6
WHEN 2=>c<="11011111";seg<="0110000";--1
WHEN 3=>c<="11101111";seg<="1101101";--2
WHEN 4=>c<="11110111";seg<="1111110";--8
WHEN 5=>c<="11111011";seg<="0110001";---
WHEN 6=>c<="11111101";seg<="1101101";--2
WHEN 7=>c<="11111110";seg<="0110000";--7
WHEN OTHERS=>c<="11111111";seg<="0000000";
END case;
END PROCESS;
END A;
