LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY yusanma IS
	PORT(
	SW:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	B:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END;
ARCHITECTURE A OF yusanma IS
BEGIN
PROCESS(SW)
BEGIN
IF SW<1001 THEN  B<=SW+"0011";
ELSE B<="0000";
END IF;
END PROCESS;
END;