LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


ENTITY lxx IS
	PORT(
		CLEAR,CLKIN:IN STD_LOGIC;
		NUM:OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		CAT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END lxx;


ARCHITECTURE BEHAVE OF lxx IS
	SIGNAL STATE:INTEGER RANGE 0 TO 8;
	BEGIN
	PROCESS(CLEAR,CLKIN)
	BEGIN
	IF CLEAR='0'THEN 
		STATE<=0;
	ELSIF (CLKIN'EVENT AND CLKIN='1')THEN
		IF STATE =8 THEN 
			STATE<=1;
		ELSE 
			STATE<=STATE+1;
		END IF;
	END IF;
END PROCESS;


PROCESS(STATE)
BEGIN
CASE STATE IS
WHEN 1=> NUM<="0110000";CAT<="01111111";--1
WHEN 2=> NUM<="1011111";CAT<="10111111";--6
WHEN 3=> NUM<="0110000";CAT<="11011111";--1
WHEN 4=> NUM<="1101101";CAT<="11101111";--2
WHEN 5=> NUM<="1111111";CAT<="11110111";--8
WHEN 6=> NUM<="0000001";CAT<="11111011";-- -
WHEN 7=> NUM<="0110000";CAT<="11111101";--1
WHEN 8=> NUM<="1011111";CAT<="11111110";--6
WHEN OTHERS=> NUM<="0000000";CAT<="00000000";
END CASE;
END PROCESS;
END BEHAVE;